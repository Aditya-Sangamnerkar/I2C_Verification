class i2cmb_coverage extends ncsu_component;

endclass : i2cmb_coverage