typedef  bit   i2c_op_t;